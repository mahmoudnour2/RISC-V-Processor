`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/25/2023 09:37:05 PM
// Design Name: 
// Module Name: memory
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module memory(input clk, input MemRead, input MemWrite,
 input [8:0] addr, input [31:0] data_in, output reg[31:0] data_out, input [2:0]func3
 );
reg [7:0] mem [511:0];
wire [8:0]offset;
assign offset = 256;



integer i;
// initial begin
 
// for(i = 0; i<512; i=i+1) begin
// mem[i] = 8'd0;
// end
 
//    {mem[256 +3],mem[256 + 2],mem[256 + 1],mem[256 + 0]} = 32'd17;
//    {mem[256 +7],mem[256 + 6],mem[256 + 5],mem[256 + 4]}  = 32'd9;
//  {mem[256 +11],mem[256 + 10],mem[256 + 9],mem[256 + 8]}  = 32'd25;
// //{mem[offset +15],mem[offset + 14],mem[offset + 13],mem[offset + 12]}  = 32'h80000000;
 
 
 
//    {mem[3],mem[2],mem[1],mem[0]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//    {mem[7],mem[6],mem[5],mem[4]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//    {mem[11],mem[10],mem[9],mem[8]} =32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//    {mem[15],mem[14],mem[13],mem[12]} =32'b000000000000_00000_010_00001_0000011 ; //lw x1, 0(x0)
//    {mem[19],mem[18],mem[17],mem[16]} =32'b000000000100_00000_010_00010_0000011 ; //lw x2, 4(x0)
//    {mem[23],mem[22],mem[21],mem[20]} =32'b000000001000_00000_010_00011_0000011 ; //lw x3, 8(x0)
//    {mem[27],mem[26],mem[25],mem[24]} =32'b0000000_00010_00001_110_00100_0110011 ; //or x4, x1, x2
//    {mem[31],mem[30],mem[29],mem[28]} =32'h00320463; //beq x4, x3, 8
//    {mem[35],mem[34],mem[33],mem[32]} =32'b0000000_00010_00001_000_00011_0110011 ; //add x3, x1, x2
//    {mem[39],mem[38],mem[37],mem[36]} =32'b0000000_00010_00011_000_00101_0110011 ; //add x5, x3, x2
//    {mem[43],mem[42],mem[41],mem[40]} =32'b0000000_00101_00000_010_01100_0100011; //sw x5, 12(x0)
//    {mem[47],mem[46],mem[45],mem[44]} =32'b000000001100_00000_010_00110_0000011 ; //lw x6, 12(x0)
//    {mem[51],mem[50],mem[49],mem[48]} =32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//    {mem[55],mem[54],mem[53],mem[52]} =32'b0000000_00001_00110_111_00111_0110011 ; //and x7, x6, x1
//    {mem[59],mem[58],mem[57],mem[56]} =32'b0100000_00010_00001_000_01000_0110011 ; //sub x8, x1, x2
//    {mem[63],mem[62],mem[61],mem[60]} =32'b0000000_00010_00001_000_00000_0110011 ; //add x0, x1, x2
//    {mem[67],mem[66],mem[65],mem[64]} =32'b0000000_00001_00000_000_01001_0110011 ; //add x9, x0, x1              
                  
                  
//         {mem[3], mem[2], mem[1], mem[0]}=32'b00000000000000001001010100010111; // auipc x10, 9
//         {mem[7], mem[6], mem[5], mem[4]}=32'b00000000000000001001010010110111; // lui x9, 9
//         {mem[11], mem[10], mem[9], mem[8]}=32'b00000000010001010000010110010011; // addi x11, x10, 4
//         {mem[15], mem[14], mem[13], mem[12]}=32'b00000000000001010000011000110011; //add x12, x10, x0
//         {mem[19], mem[18], mem[17], mem[16]}=32'b00000000100000000000000011101111; //jal ra,8
//         {mem[23], mem[22], mem[21], mem[20]}=32'b00000000000100000000000001110011; // ebreak
//         {mem[27], mem[26], mem[25], mem[24]}=32'b00001000101101010000110001100011; //beq x10, x11, 152
//         {mem[31], mem[30], mem[29], mem[28]}=32'b00000000101101010001010001100011 ;//bne x10, x11, 8
//         {mem[35], mem[34], mem[33], mem[32]}=32'b00000000000000000000000001110011; // ecall
//         {mem[39], mem[38], mem[37], mem[36]}=32'b00000011001000000000001100010011; //addi x6, x0, 50
//         {mem[43], mem[42], mem[41], mem[40]}=32'b00000000001000110001001100010011; //slli x6, x6, 2
//         {mem[47], mem[46], mem[45], mem[44]}=32'b00000000001000000000001110010011 ; //addi x7, x0, 2
//         {mem[51], mem[50], mem[49], mem[48]}=32'b00000000011100000000000000100011;//sb x7, 0(x0)
//         {mem[55], mem[54], mem[53], mem[52]}=32'b00000000101000000001000000100011; //sh x10, 0(x0)
//         {mem[59], mem[58], mem[57], mem[56]}=32'b00000000101000000010000000100011; // sw x10, 0(x0)
//         {mem[63], mem[62], mem[61], mem[60]}=32'b00000000000000000000111000000011; // lb x28, 0(x0)
//         {mem[67], mem[66], mem[65], mem[64]}=32'b00000000000000000001111010000011;//lh x29, 0(x0)
//         {mem[71], mem[70], mem[69], mem[68]}=32'b00000000000000000010111100000011; //lw x30, 0(x0)
//         {mem[75], mem[74], mem[73], mem[72]}=32'b00000000000000000100111110000011; //lbu x31, 0(x0)
//         {mem[79], mem[78], mem[77], mem[76]}=32'b00000000000000000101001100000011; //lhu x6, 0(x0)
//         {mem[83], mem[82], mem[81], mem[80]}=32'b00000110101101100101000001100011; // bge x12, x11, 96
//         {mem[87], mem[86], mem[85], mem[84]}=32'b00000100110001011100111001100011; //blt x11, x12, 92
//         {mem[91], mem[90], mem[89], mem[88]}=32'b00000100101101100111110001100011; //bgeu x12, x11, 88
//         {mem[95], mem[94], mem[93], mem[92]}=32'b00000100110001011110101001100011; //bltu x11, x12, 84
//         {mem[99], mem[98], mem[97], mem[96]}=32'b11111001110001100011001100010011; //sltiu x6, x12, -100
//         {mem[103], mem[102], mem[101], mem[100]}=32'b00000000001100110100111000010011; //xori x28, x6, 3
//         {mem[107], mem[106], mem[105], mem[104]}=32'b00000000010111100110111000010011; //ori x28, x28, 5
//         {mem[111], mem[110], mem[109], mem[108]}=32'b00000000010111100111111000010011; //andi x28, x28, 5
//         {mem[115], mem[114], mem[113], mem[112]}=32'b00000000000111100101111000010011; //srli x28, x28, 1
//         {mem[119], mem[118], mem[117], mem[116]}=32'b00000010100011100000111000010011; //addi x28, x28, 40
//         {mem[123], mem[122], mem[121], mem[120]}=32'b01000000001011100101111000010011; //srai x28, x28, 2
//         {mem[127], mem[126], mem[125], mem[124]}=32'b00000000001100000000001110010011; //addi x7, x0, 3
//         {mem[131], mem[130], mem[129], mem[128]}=32'b01000000011111100000111000110011; // sub x28, x28, x7
//         {mem[135], mem[134], mem[133], mem[132]}=32'b00000001110011100001111000110011; //sll x28, x28, x28
//         {mem[139], mem[138], mem[137], mem[136]}=32'b00000001110011100010111100110011; //slt x30, x28, x28
//         {mem[143], mem[142], mem[141], mem[140]}=32'b00000000011000000000111010010011; //addi x29, x0, 6
//         {mem[147], mem[146], mem[145], mem[144]}=32'b00000001110011101011111100110011; //sltu x30, x29, x28
//         {mem[151], mem[150], mem[149], mem[148]}=32'b00000001110111110100111100110011; //xor x30, x30, x29
//         {mem[155], mem[154], mem[153], mem[152]}=32'b00000000010011110001111100010011; //slli x30, x30, 4
//         {mem[159], mem[158], mem[157], mem[156]}=32'b00000000011111110101111100110011; //srl x30, x30, x7
//         {mem[163], mem[162], mem[161], mem[160]}=32'b01000000011111110101111100110011; //sra x30, x30, x7
//         {mem[167], mem[166], mem[165], mem[164]}=32'b00000000011111110110111100110011; //or x30, x30, x7
//         {mem[171], mem[170], mem[169], mem[168]}=32'b00000001110111110111111100110011; //and x30, x30, x29
//         {mem[175], mem[174], mem[173], mem[172]}=32'b00000000000000000000000000001111;// fence
//         {mem[179], mem[178], mem[177], mem[176]}=32'b00000000000000001000000001100111; // jalr x0, 0(x1)
                  
//end    


//store
 always @(negedge clk) begin
 if(MemWrite ==1) begin
    case(func3)
    3'b000: mem[256 +addr] = data_in[7:0];//SB
    3'b001: begin mem[256 +addr] = data_in[7:0];
    mem[256 +addr+1]= data_in[15:8];//SH
    end
    3'b010: begin mem[256 + addr] = data_in[7:0];
    mem[256 + addr + 1]=data_in[15:8]; 
    mem[256 + addr + 2]=data_in[23:16];
    mem[256 + addr + 3]=data_in[31:24];
    end //SW
    endcase
 end
 end

 
 always @(*) begin
 if(!clk) begin
     if(MemRead == 1)begin
        case(func3)
        //3'b000: data_out  <=  {{24{mem[addr][7]}},mem[addr]};//LB
        3'b000: data_out  <=  {(mem[256 +addr][7]==1'b1)?24'hffffff:24'h000000,mem[256 +addr]};//LB
        //3'b001: data_out  <=  {{16{mem[addr][15]}},mem[addr+1],mem[addr]};//LH
        3'b001: data_out  <=  {(mem[256 +addr+1][7]==1'b1)?16'hffff:16'h0000,mem[256 +addr+1],mem[offset +addr]};//LH
        3'b010: begin
            data_out  <=  {mem[256 +addr+3],mem[256 +addr+2],mem[256 +addr+1],mem[256 +addr]};//LW
        end
        3'b100: data_out  <=  {24'd0,mem[256 +addr]};//LBU
        3'b101: data_out  <=  {16'd0,mem[256 +addr+1],mem[256 +addr]};//LHU
        endcase
     end
  end
  else data_out <= {mem[addr+3],mem[addr+2],mem[addr+1],mem[addr]};
 end
 
 
 initial begin                    
                       
 for(i = 0; i<512; i=i+1) begin   
 mem[i] = 8'd0;                   
 end              
                                                                                                                                                                                      
 {mem[3], mem[2], mem[1], mem[0]} = 32'h01663c33; // sltu x24, x12, x22                            
 {mem[7], mem[6], mem[5], mem[4]} = 32'h0055a233; // slt x4, x11, x5                               
 {mem[11], mem[10], mem[9], mem[8]} = 32'hb094e717; // auipc x14, 723278                           
 {mem[15], mem[14], mem[13], mem[12]} = 32'hc83894b7; // lui x9, 820105                            
 {mem[19], mem[18], mem[17], mem[16]} = 32'h005b5c93; // srli x25, x22, 1252                       
 {mem[23], mem[22], mem[21], mem[20]} = 32'hfb07cb83; // lbu x23, -80(x15)                         
 {mem[27], mem[26], mem[25], mem[24]} = 32'h01592e33; // slt x28, x18, x21                         
 {mem[31], mem[30], mem[29], mem[28]} = 32'hb605d183; // lhu x3, -1184(x11)                        
 {mem[35], mem[34], mem[33], mem[32]} = 32'h098cd983; // lhu x19, 152(x25)                         
 {mem[39], mem[38], mem[37], mem[36]} = 32'h007bc863; // blt x23, x7, 1056                         
 {mem[43], mem[42], mem[41], mem[40]} = 32'h418a8f93; // addi x31, x21, 1048                       
 {mem[47], mem[46], mem[45], mem[44]} = 32'h6ce31a63; // bne x6, x14, 1748                         
 {mem[51], mem[50], mem[49], mem[48]} = 32'h01c4b833; // sltu x16, x9, x28                         
 {mem[55], mem[54], mem[53], mem[52]} = 32'h150008ef; // add x31, x11, x19                         
 {mem[59], mem[58], mem[57], mem[56]} = 32'h0077fbb3; // jal x17, 336                              
 {mem[63], mem[62], mem[61], mem[60]} = 32'h36d4ce63; // and x23, x15, x7                          
 {mem[67], mem[66], mem[65], mem[64]} = 32'hcdd35097; // blt x9, x13, 892                          
 {mem[71], mem[70], mem[69], mem[68]} = 32'h009b5c13; // auipc x1, 843061                          
 {mem[75], mem[74], mem[73], mem[72]} = 32'h6e964263; // srli x24, x22, -57                        
 {mem[79], mem[78], mem[77], mem[76]} = 32'h36c11623; // blt x12, x9, 1764                         
 {mem[83], mem[82], mem[81], mem[80]} = 32'h004482b3; // add x5, x9, x4                            
 {mem[87], mem[86], mem[85], mem[84]} = 32'h00879693; // slli x13, x15, -1611                      
 {mem[91], mem[90], mem[89], mem[88]} = 32'h15d70837; // lui x16, 89456                            
 {mem[95], mem[94], mem[93], mem[92]} = 32'h01966fb3; // or x31, x12, x25                          
 {mem[99], mem[98], mem[97], mem[96]} = 32'h36c11623; // sh x12, 876(x2)                           
 {mem[103], mem[102], mem[101], mem[100]} = 32'h748003ef; // jal x7, 1864                          
 {mem[107], mem[106], mem[105], mem[104]} = 32'hc3780993; // addi x19, x16, -969                   
 {mem[111], mem[110], mem[109], mem[108]} = 32'h7907d7b7; // lui x15, 495741                       
 {mem[115], mem[114], mem[113], mem[112]} = 32'hcf341823; // sh x19, -784(x8)                      
 {mem[119], mem[118], mem[117], mem[116]} = 32'h25c00ee7; // jalr x29, 604                         


// {mem[3], mem[2], mem[1], mem[0]} =32'b0000000_00000_00000_000_00000_0110011;// noop   
// {mem[7], mem[6], mem[5], mem[4]} = 32'hffb00113; // Addi x2,x0,-5 
// {mem[11], mem[10], mem[9], mem[8]}=32'h00400493; // Addi x9,x0,4  
// {mem[15], mem[14], mem[13], mem[12]}=  32'h00302223; // Sw x3,4(x0)      
// {mem[19], mem[18], mem[17], mem[16]} = 32'h00200023; // Sb x2, 0(x0)     
// {mem[23], mem[22], mem[21], mem[20]} = 32'h00000203;//Lb x4, 0(x0)       
// {mem[27], mem[26], mem[25], mem[24]} = 32'h00201283;// Lh x5, 2(x0)      
// {mem[31], mem[30], mem[29], mem[28]} = 32'h00402303; //Lw x6, 4(x0)      
// {mem[35], mem[34], mem[33], mem[32]} = 32'h00855463; //Bge x10,x8,8        
// {mem[39], mem[38], mem[37], mem[36]} = 32'h00a12213; // Slti x4,x2,10         
// {mem[43], mem[42], mem[41], mem[40]} = 32'hff613213; // Sltiu x4, x2,-10   
// {mem[47], mem[46], mem[45], mem[44]} = 32'h01024213; // Xori x4,x4,16      
// {mem[51], mem[50], mem[49], mem[48]} = 32'h01b4e313; // Ori x6,x9, 27                                         
// {mem[55], mem[54], mem[53], mem[52]} = 32'h000df393; // Andi x7,x27,0                                         
// {mem[59], mem[58], mem[57], mem[56]} = 32'h40a4d913; // Srai x18,x9,10                                            
// {mem[63], mem[62], mem[61], mem[60]} = 32'h40950433; // Sub x8,x10,x9    
// {mem[67], mem[66], mem[65], mem[64]} = 32'h00481d33; //Sll x26,x16,x4    
// {mem[71], mem[70], mem[69], mem[68]} = 32'h02a50463; // Beq x10,x10, 40  
// {mem[75], mem[74], mem[73], mem[72]} = 32'h0042c533; // Xor x10,x5,x4    
// {mem[79], mem[78], mem[77], mem[76]} =  32'h0031d1b3; // Srl x3,x3,x3                                         
// {mem[83], mem[82], mem[81], mem[80]} =  32'h0090e263; //Bltu x1,x9,4     
// {mem[87], mem[86], mem[85], mem[84]}=  32'h40215133; // Sra x2,x2,x2     
// {mem[91], mem[90], mem[89], mem[88]}= 32'h0041e1b3; // Or x3,x3,x4  
// {mem[95], mem[94], mem[93], mem[92]}=  32'b00000000000100000000000001110011;// ebreak 




end



endmodule
































































